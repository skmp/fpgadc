localparam REG0_BANK0   = 6'd0;
localparam REG1_BANK0   = 6'd1;
localparam REG2_BANK0   = 6'd2;
localparam REG3_BANK0   = 6'd3;
localparam REG4_BANK0   = 6'd4;
localparam REG5_BANK0   = 6'd5;
localparam REG6_BANK0   = 6'd6;
localparam REG7_BANK0   = 6'd7;
localparam REG8         = 6'd8;
localparam REG9         = 6'd9;
localparam REG10        = 6'd10;
localparam REG11        = 6'd11;
localparam REG12        = 6'd12;
localparam REG13        = 6'd13;
localparam REG14        = 6'd14;
localparam REG15        = 6'd15;

localparam REG0_BANK1   = 6'd16;
localparam REG1_BANK1   = 6'd17;
localparam REG2_BANK1   = 6'd18;
localparam REG3_BANK1   = 6'd19;
localparam REG4_BANK1   = 6'd20;
localparam REG5_BANK1   = 6'd21;
localparam REG6_BANK1   = 6'd21;
localparam REG7_BANK1   = 6'd23;

localparam REG_MACL     = 6'd24;
localparam REG_MACH     = 6'd25;

localparam REG_FPUL     = 6'd26;

localparam REG_CONST_0  = 6'd31;
localparam REG_CONST_1  = 6'd32;

localparam REG_FR0      = 6'd32;
localparam REG_FR1      = 6'd33;
localparam REG_FR2      = 6'd34;
localparam REG_FR3      = 6'd35;
localparam REG_FR4      = 6'd36;
localparam REG_FR5      = 6'd37;
localparam REG_FR6      = 6'd38;
localparam REG_FR7      = 6'd39;
localparam REG_FR8      = 6'd40;
localparam REG_FR9      = 6'd41;
localparam REG_FR10     = 6'd42;
localparam REG_FR11     = 6'd43;
localparam REG_FR12     = 6'd44;
localparam REG_FR13     = 6'd45;
localparam REG_FR14     = 6'd46;
localparam REG_FR15     = 6'd47;

localparam REG_XFR0     = 6'd48;
localparam REG_XFR1     = 6'd49;
localparam REG_XFR2     = 6'd50;
localparam REG_XFR3     = 6'd51;
localparam REG_XFR4     = 6'd52;
localparam REG_XFR5     = 6'd53;
localparam REG_XFR6     = 6'd54;
localparam REG_XFR7     = 6'd55;
localparam REG_XFR8     = 6'd56;
localparam REG_XFR9     = 6'd57;
localparam REG_XFR10    = 6'd58;
localparam REG_XFR11    = 6'd59;
localparam REG_XFR12    = 6'd60;
localparam REG_XFR13    = 6'd61;
localparam REG_XFR14    = 6'd62;
localparam REG_XFR15    = 6'd63;
