localparam ADD = 6'd0;
localparam SUBTRACT = 6'd1;
localparam MULTIPLY = 6'd2;
localparam DIVIDE = 6'd3;

localparam AND = 6'd4;
localparam OR = 6'd5;
localparam XOR = 6'd6;

localparam LOAD8 = 6'd8;
localparam STORE8 = 6'd9;
localparam LOAD16 = 6'd10;
localparam STORE16 = 6'd11;
localparam LOAD32 = 6'd12;
localparam STORE32 = 6'd13;

localparam ILLEGAL = 6'd63;
